
// GPIO port width
//  min value 1
//  max value 32
`define SM_GPIO_WIDTH       4

